/*************************************************************************
	> File Name: IFU.v
	> Author: Jensen
	> Mail: 1624839259@qq.com 
	> Created Time: 2024年10月06日 星期日 16时04分06秒
 ************************************************************************/
module ysyx_24090018_IFU #(ADDR_WIDTH = 32, DATA_WIDTH = 32)(
  input clk,
  input [ADDR_WIDTH-1 : 0] pc,
  output [DATA_WIDTH-1 : 0] inst_o
);


endmodule
