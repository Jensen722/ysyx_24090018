/*************************************************************************
	> File Name: add_32bit.v
	> Author: Jensen
	> Mail: 1624839259@qq.com 
	> Created Time: 2024年12月06日 星期五 19时27分33秒
 ************************************************************************/
module add_32bit(
  input [31:0] a,
  input [31:0] b,
  output [31:0] s
);
  wire carry;
  assign {carry, s} = a + b;  //先设计成串行进位加法器，后面再更改加法器位进位选择加法
  //器，减少延时
  //不考虑进位，也不考虑溢出

endmodule
